
module ece120_not(
    input logic op,
    output logic res
    );
    assign res = ~op;
endmodule